`timescale 1ns / 1ps


module reverse_circuit(

    );
endmodule
